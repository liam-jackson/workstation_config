
bindkey -R " "-"~" self-insert
bindkey -R "\M-^@"-"\M-^?" self-insert
bindkey "^_" undo
bindkey "^?" backward-delete-char
bindkey "^[ " expand-history
bindkey "^[_" insert-last-word
bindkey "^[-" neg-argument
bindkey "^[," _history-complete-newer
bindkey "^[!" expand-history
bindkey "^[?" which-command
bindkey "^[." insert-last-word
bindkey "^['" quote-line
bindkey "^[[0n" reset-prompt
bindkey "^[[2~" overwrite-mode
bindkey "^[[200~" bracketed-paste
bindkey "^[[3~" delete-char
bindkey "^[[A" up-line-or-history
bindkey "^[[B" down-line-or-history
bindkey "^[[C" forward-char
bindkey "^[[D" backward-char
bindkey "^[/" _history-complete-older
bindkey "^[\"" quote-region
bindkey "^[\$" spell-word
bindkey "^[^_" copy-prev-word
bindkey "^[^?" backward-kill-word
bindkey "^[^D" list-choices
bindkey "^[^G" send-break
bindkey "^[^H" backward-kill-word
bindkey "^[^I" self-insert-unmeta
bindkey "^[^J" self-insert-unmeta
bindkey "^[^L" clear-screen
bindkey "^[^M" self-insert-unmeta
bindkey "^[<" beginning-of-buffer-or-history
bindkey "^[>" end-of-buffer-or-history
bindkey "^[|" vi-goto-column
bindkey "^[~" _bash_complete-word
bindkey "^[0" digit-argument
bindkey "^[1" digit-argument
bindkey "^[2" digit-argument
bindkey "^[3;5~" delete-char
bindkey "^[3" digit-argument
bindkey "^[4" digit-argument
bindkey "^[5" digit-argument
bindkey "^[6" digit-argument
bindkey "^[7" digit-argument
bindkey "^[8" digit-argument
bindkey "^[9" digit-argument
bindkey "^[a" accept-and-hold
bindkey "^[A" accept-and-hold
bindkey "^[b" backward-word
bindkey "^[B" backward-word
bindkey "^[C" capitalize-word
bindkey "^[c" fzf-cd-widget
bindkey "^[d" kill-word
bindkey "^[D" kill-word
bindkey "^[f" forward-word
bindkey "^[F" forward-word
bindkey "^[g" get-line
bindkey "^[G" get-line
bindkey "^[ga" fzf-git-add-files
bindkey "^[h" run-help
bindkey "^[H" run-help
bindkey "^[l" down-case-word
bindkey "^[L" down-case-word
bindkey "^[n" history-search-forward
bindkey "^[N" history-search-forward
bindkey "^[OA" up-line-or-history
bindkey "^[OB" down-line-or-history
bindkey "^[OC" forward-char
bindkey "^[OD" backward-char
bindkey "^[OF" end-of-line
bindkey "^[OH" beginning-of-line
bindkey "^[p" history-search-backward
bindkey "^[P" history-search-backward
bindkey "^[q" push-line
bindkey "^[Q" push-line
bindkey "^[s" spell-word
bindkey "^[S" spell-word
bindkey "^[t" transpose-words
bindkey "^[T" transpose-words
bindkey "^[u" up-case-word
bindkey "^[U" up-case-word
bindkey "^[w" copy-region-as-kill
bindkey "^[W" copy-region-as-kill
bindkey "^[x" execute-named-cmd
bindkey "^[y" yank-pop
bindkey "^[z" execute-last-named-cmd
bindkey "^@" set-mark-command
bindkey "^\\\\" fzf-select-widget
bindkey "^A" beginning-of-line
bindkey "^B" backward-char
bindkey "^D" delete-char-or-list
bindkey "^E" end-of-line
bindkey "^F" forward-char
bindkey "^G" send-break
bindkey "^G^B" fzf-git-branches-widget
bindkey "^G^E" fzf-git-each_ref-widget
bindkey "^G^F" fzf-git-files-widget
bindkey "^G^H" fzf-git-hashes-widget
bindkey "^G^L" fzf-git-lreflogs-widget
bindkey "^G^R" fzf-git-remotes-widget
bindkey "^G^S" fzf-git-stashes-widget
bindkey "^G^T" fzf-git-tags-widget
bindkey "^Gb" fzf-git-branches-widget
bindkey "^Ge" fzf-git-each_ref-widget
bindkey "^Gf" fzf-git-files-widget
bindkey "^Gh" fzf-git-hashes-widget
bindkey "^Gl" fzf-git-lreflogs-widget
bindkey "^Gr" fzf-git-remotes-widget
bindkey "^Gs" fzf-git-stashes-widget
bindkey "^Gt" fzf-git-tags-widget
bindkey "^H" fzf-man-widget
bindkey "^I" fzf-tab-complete
bindkey "^J" accept-line
bindkey "^K" kill-line
bindkey "^L" clear-screen
bindkey "^M" accept-line
bindkey "^N" down-line-or-history
bindkey "^O" accept-line-and-down-history
bindkey "^P" up-line-or-history
bindkey "^Q" push-line
bindkey "^R" fzf-history-widget
bindkey "^S" history-incremental-search-forward
bindkey "^T" fzf-file-widget
bindkey "^U" kill-whole-line
bindkey "^V" quoted-insert
bindkey "^W" backward-kill-word
bindkey "^X?" _complete_debug
bindkey "^X." fzf-tab-debug
bindkey "^X*" expand-word
bindkey "^X^B" vi-match-bracket
bindkey "^X^F" vi-find-next-char
bindkey "^X^J" vi-join
bindkey "^X^K" kill-buffer
bindkey "^X^N" infer-next-history
bindkey "^X^O" overwrite-mode
bindkey "^X^R" _read_comp
bindkey "^X^U" undo
bindkey "^X^V" vi-cmd-mode
bindkey "^X^X" exchange-point-and-mark
bindkey "^X=" what-cursor-position
bindkey "^X~" _bash_list-choices
bindkey "^Xa" _expand_alias
bindkey "^XC" _correct_filename
bindkey "^Xc" _correct_word
bindkey "^Xd" _list_expansions
bindkey "^Xe" _expand_word
bindkey "^Xg" list-expand
bindkey "^XG" list-expand
bindkey "^Xh" _complete_help
bindkey "^Xm" _most_recent_file
bindkey "^Xn" _next_tags
bindkey "^Xr" history-incremental-search-backward
bindkey "^Xs" history-incremental-search-forward
bindkey "^Xt" _complete_tag
bindkey "^Xu" undo
bindkey "^Y" yank
