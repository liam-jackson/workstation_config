bindkey "^[\$" spell-word
bindkey "^[0" digit-argument
bindkey "^[[0n" reset-prompt
bindkey "^[1" digit-argument
bindkey "^[[200~" bracketed-paste
bindkey "^[2" digit-argument
bindkey "^[[2~" overwrite-mode
bindkey "^[3;5~" delete-char
bindkey "^[[3~" delete-char
bindkey "^[3" digit-argument
bindkey "^[4" digit-argument
bindkey "^[5" digit-argument
bindkey "^[6" digit-argument
bindkey "^[7" digit-argument
bindkey "^[8" digit-argument
bindkey "^[9" digit-argument
bindkey "^[a" accept-and-hold
bindkey "^[A" accept-and-hold
bindkey "^A" beginning-of-line
bindkey "^[[A" up-line-or-history
bindkey "^?" backward-delete-char
bindkey "^[^?" backward-kill-word
bindkey "^[~" _bash_complete-word
bindkey "^B" backward-char
bindkey "^[b" backward-word
bindkey "^[B" backward-word
bindkey "^[[B" down-line-or-history
bindkey "^[<" beginning-of-buffer-or-history
bindkey "^[C" capitalize-word
bindkey "^[[C" forward-char
bindkey "^[c" fzf-cd-widget
bindkey "^[^_" copy-prev-word
bindkey "^[[D" backward-char
bindkey "^D" delete-char-or-list
bindkey "^[d" kill-word
bindkey "^[D" kill-word
bindkey "^[^D" list-choices
bindkey "^E" end-of-line
bindkey "^[>" end-of-buffer-or-history
bindkey "^[ " expand-history
bindkey "^[!" expand-history
bindkey "^F" forward-char
bindkey "^[f" forward-word
bindkey "^[F" forward-word
bindkey "^\\\\" fzf-select-widget
bindkey "^[ga" fzf-git-add-files
bindkey "^Gb" fzf-git-branches-widget
bindkey "^G^B" fzf-git-branches-widget
bindkey "^Ge" fzf-git-each_ref-widget
bindkey "^G^E" fzf-git-each_ref-widget
bindkey "^Gf" fzf-git-files-widget
bindkey "^G^F" fzf-git-files-widget
bindkey "^[g" get-line
bindkey "^[G" get-line
bindkey "^Gh" fzf-git-hashes-widget
bindkey "^G^H" fzf-git-hashes-widget
bindkey "^Gl" fzf-git-lreflogs-widget
bindkey "^G^L" fzf-git-lreflogs-widget
bindkey "^Gr" fzf-git-remotes-widget
bindkey "^G^R" fzf-git-remotes-widget
bindkey "^[^G" send-break
bindkey "^G" send-break
bindkey "^Gs" fzf-git-stashes-widget
bindkey "^G^S" fzf-git-stashes-widget
bindkey "^Gt" fzf-git-tags-widget
bindkey "^G^T" fzf-git-tags-widget
bindkey "^[^H" backward-kill-word
bindkey "^H" fzf-man-widget
bindkey "^[," _history-complete-newer
bindkey "^[/" _history-complete-older
bindkey "^[h" run-help
bindkey "^[H" run-help
bindkey "^I" fzf-tab-complete
bindkey "^[." insert-last-word
bindkey "^[_" insert-last-word
bindkey "^[^I" self-insert-unmeta
bindkey "^J" accept-line
bindkey "^[^J" self-insert-unmeta
bindkey "^K" kill-line
bindkey "^[^L" clear-screen
bindkey "^L" clear-screen
bindkey "^[l" down-case-word
bindkey "^[L" down-case-word
bindkey "^M" accept-line
bindkey "^[^M" self-insert-unmeta
bindkey "^N" down-line-or-history
bindkey "^[-" neg-argument
bindkey "^[n" history-search-forward
bindkey "^[N" history-search-forward
bindkey "^O" accept-line-and-down-history
bindkey "^[OA" up-line-or-history
bindkey "^[OB" down-line-or-history
bindkey "^[OC" forward-char
bindkey "^[OD" backward-char
bindkey "^[OF" end-of-line
bindkey "^[OH" beginning-of-line
bindkey "^[p" history-search-backward
bindkey "^[P" history-search-backward
bindkey "^P" up-line-or-history
bindkey "^[q" push-line
bindkey "^[Q" push-line
bindkey "^Q" push-line
bindkey "^['" quote-line
bindkey "^[\"" quote-region
bindkey "^R" fzf-history-widget
bindkey -R "\M-^@"-"\M-^?" self-insert
bindkey -R " "-"~" self-insert
bindkey "^@" set-mark-command
bindkey "^S" history-incremental-search-forward
bindkey "^[s" spell-word
bindkey "^[S" spell-word
bindkey "^T" fzf-file-widget
bindkey "^[t" transpose-words
bindkey "^[T" transpose-words
bindkey "^U" kill-whole-line
bindkey "^_" undo
bindkey "^[u" up-case-word
bindkey "^[U" up-case-word
bindkey "^[|" vi-goto-column
bindkey "^V" quoted-insert
bindkey "^W" backward-kill-word
bindkey "^[w" copy-region-as-kill
bindkey "^[W" copy-region-as-kill
bindkey "^[?" which-command
bindkey "^Xa" _expand_alias
bindkey "^X~" _bash_list-choices
bindkey "^X^B" vi-match-bracket
bindkey "^XC" _correct_filename
bindkey "^Xc" _correct_word
bindkey "^X?" _complete_debug
bindkey "^Xd" _list_expansions
bindkey "^Xe" _expand_word
bindkey "^[x" execute-named-cmd
bindkey "^X*" expand-word
bindkey "^X^F" vi-find-next-char
bindkey "^X." fzf-tab-debug
bindkey "^Xg" list-expand
bindkey "^XG" list-expand
bindkey "^Xh" _complete_help
bindkey "^X^J" vi-join
bindkey "^X^K" kill-buffer
bindkey "^Xm" _most_recent_file
bindkey "^X^N" infer-next-history
bindkey "^Xn" _next_tags
bindkey "^X^O" overwrite-mode
bindkey "^Xr" history-incremental-search-backward
bindkey "^X^R" _read_comp
bindkey "^Xs" history-incremental-search-forward
bindkey "^Xt" _complete_tag
bindkey "^Xu" undo
bindkey "^X^U" undo
bindkey "^X^V" vi-cmd-mode
bindkey "^X=" what-cursor-position
bindkey "^X^X" exchange-point-and-mark
bindkey "^Y" yank
bindkey "^[y" yank-pop
bindkey "^[z" execute-last-named-cmd
